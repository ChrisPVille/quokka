module cpu_control(
    input clk,
    input rst_n,
    input[15:0] A,
    input[7:0] D
    );

    always@(posedge clk or negedge rst_n) begin
        
    end

endmodule
