module top(
    );


endmodule
